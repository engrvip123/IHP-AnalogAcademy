* Extracted by KLayout with SG13G2 LVS runset on : 13/02/2025 13:18

.SUBCKT two_stage_OTA_layout vss vdd dn3 iout vout dn2 v+ v\x2d vss$1 dn4
M$1 vss dn3 dn3 vss sg13_lv_nmos L=9.75u W=0.72u AS=0.2448p AD=0.2448p PS=2.12u
+ PD=2.12u
M$2 vss dn3 dn4 vss sg13_lv_nmos L=9.75u W=0.72u AS=0.2448p AD=0.2448p PS=2.12u
+ PD=2.12u
M$3 vss$1 dn4 vout vss sg13_lv_nmos L=9.75u W=28.8u AS=6.552p AD=6.552p
+ PS=37.82u PD=37.82u
M$7 vdd iout iout \$3 sg13_lv_pmos L=2.08u W=75u AS=15.65625p AD=15.65625p
+ PS=87.715u PD=87.715u
M$15 vdd iout vout \$3 sg13_lv_pmos L=2.08u W=75u AS=15.65625p AD=15.65625p
+ PS=87.715u PD=87.715u
M$23 vdd vdd dn2 \$2 sg13_lv_pmos L=3.7u W=14.56u AS=4.9504p AD=4.9504p
+ PS=31.84u PD=31.84u
M$25 dn2 v+ dn4 \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p PS=15.92u
+ PD=15.92u
M$26 dn2 v\x2d dn3 \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$27 dn4 vdd vdd \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$28 dn3 vdd vdd \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$35 dn2 iout vdd \$38 sg13_lv_pmos L=1.95u W=5.3u AS=1.802p AD=1.802p
+ PS=11.28u PD=11.28u
C$36 \$7 vout cap_cmim w=22.295u l=22.295u A=497.067025p P=89.18u m=1
R$37 \$3 vdd ntap1 A=27.435p P=177u
R$38 \$2 vdd ntap1 A=28.7556p P=185.52u
R$39 \$38 vdd ntap1 A=7.5826p P=48.92u
R$40 vss vss$1 ptap1 A=25.19p P=201.52u
.ENDS two_stage_OTA_layout
