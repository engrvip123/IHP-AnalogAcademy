* Extracted by KLayout with SG13G2 LVS runset on : 13/02/2025 13:49

.SUBCKT input_stage dn3|dn4|vss vdd dn2 iout
M$1 dn3|dn4|vss dn3|dn4|vss dn3|dn4|vss \$1 sg13_lv_nmos L=9.75u W=1.44u
+ AS=0.4896p AD=0.4896p PS=4.24u PD=4.24u
M$3 dn2 iout vdd \$6 sg13_lv_pmos L=1.95u W=5.3u AS=1.802p AD=1.802p PS=11.28u
+ PD=11.28u
R$4 \$6 vdd ntap1 A=21.5031p P=43.5u
R$5 \$1 dn3|dn4|vss ptap1 A=15.54345p P=53.44u
.ENDS input_stage
