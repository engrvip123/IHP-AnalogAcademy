** sch_path: /home/pedersen/projects/IHP-AnalogAcademy/modules/module_1_bandgap_reference/part_3_layout/OTA_layout/output_stage/schematic_mod/output_stage.sch
.subckt output_stage vdd iout vout vss dn4
*.PININFO vdd:B iout:B vout:B vss:B dn4:B
M7 vout iout vdd bulk3 sg13_lv_pmos l=2.08u w=75u ng=8 m=1
M6 vout dn4 vss bulk2 sg13_lv_nmos l=9.75u w=28.8u ng=4 m=1
M9 iout iout vdd bulk3 sg13_lv_pmos l=2.08u w=75u ng=8 m=1
C2 dn4 vout cap_cmim w=22.295e-6 l=22.295e-6 m=1
R2 vss bulk2 ptap1 A = 68.4036e-12, P = 0.24264e-3
R5 vdd bulk3 ntap1 A = 95.5222e-12, P = 0.21292e-3
.ends
.end

