** sch_path: /home/pedersen/projects/IHP-AnalogAcademy/modules/module_1_bandgap_reference/part_3_layout/OTA_layout/input_pair/schematic_mod/input_common_centroid.sch
.subckt input_common_centroid v- v+ vdd dn3 dn4
*.PININFO v-:B v+:B vdd:B dn3:B dn4:B
M1 dn3 v- dn2 bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M2 dn4 v+ dn2 bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M8 dn4 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M10 dn3 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M15 dn2 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M16 dn2 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
R1 vdd bulk ntap1 A = 0.1979248e-9 P = 0.2436e-3

.ends
.end
