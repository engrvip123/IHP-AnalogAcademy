* Extracted by KLayout with SG13G2 LVS runset on : 18/03/2025 08:57

.SUBCKT input_common_centroid v+ v\x2d vdd dn4 dn3
M$1 vdd vdd \$6 \$27 sg13_lv_pmos L=3.7u W=14.56u AS=4.9504p AD=4.9504p
+ PS=31.84u PD=31.84u
M$2 \$6 v+ dn4 \$27 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p PS=15.92u
+ PD=15.92u
M$3 dn4 vdd vdd \$27 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$5 \$6 v\x2d dn3 \$27 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$6 dn3 vdd vdd \$27 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
.ENDS input_common_centroid
