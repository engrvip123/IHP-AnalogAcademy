** sch_path: /home/pedersen/projects/IHP-AnalogAcademy/modules/module_0_foundations/xschem/nmos_intrin.sch
**.subckt nmos_intrin
XM2 Vout net2 GND GND sg13_lv_nmos w=46.54 l=3.25u ng=1 m=5
I1 Vdd net1 13.96e-6
XM5 net1 net1 GND GND sg13_lv_nmos w=46.54 l=3.25u ng=1 m=5
Vdd Vdd GND 1.2
C1 Vout GND 1p m=1
Vin net1 net2 AC
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt



.control
op
ac dec 20 1 1e9
save all
let Av = db(v(vout))
write output_file.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
