* Extracted by KLayout with SG13G2 LVS runset on : 27/03/2025 16:05

.SUBCKT output_stage vout dn4 vdd iout vss vout$1 vout$2 dn4$1
M$1 vss dn4$1 vout$2 \$1 sg13_lv_nmos L=9.75u W=28.8u AS=6.552p AD=6.552p
+ PS=37.82u PD=37.82u
M$5 vdd iout iout \$4 sg13_lv_pmos L=2.08u W=75u AS=15.65625p AD=15.65625p
+ PS=87.715u PD=87.715u
M$13 vdd iout vout$1 \$4 sg13_lv_pmos L=2.08u W=75u AS=15.65625p AD=15.65625p
+ PS=87.715u PD=87.715u
C$21 dn4 vout cap_cmim w=22.295u l=22.295u A=497.067025p P=89.18u m=1
R$22 \$4 vdd ntap1 A=27.435p P=177u
R$23 \$1 vss ptap1 A=25.19p P=201.52u
.ENDS output_stage
