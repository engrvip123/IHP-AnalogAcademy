** sch_path: /home/pedersen/projects/IHP-AnalogAcademy/modules/module_1_bandgap_reference/part_1_OTA/xschem/two_stage_OTA.sch
**.subckt two_stage_OTA v- v+ itail vdd vss vdd iout vout
*.iopin v-
*.iopin v+
*.iopin itail
*.iopin vdd
*.iopin vss
*.iopin vdd
*.iopin iout
*.iopin vout
XM4 net3 net1 vss vss sg13_lv_nmos w=0.50u l=9.75u ng=1 m=1
XM3 net1 net1 vss vss sg13_lv_nmos w=0.50u l=9.75u ng=1 m=1
XM1 net1 v- net2 vdd sg13_lv_pmos w=6.96u l=3.25u ng=4 m=1
XM2 net3 v+ net2 vdd sg13_lv_pmos w=6.96u l=3.25u ng=4 m=1
XM5 net2 itail vdd vdd sg13_lv_pmos w=3u l=130n ng=1 m=1
XM8 itail itail vdd vdd sg13_lv_pmos w=3u l=130n ng=1 m=1
XM7 vout bias vdd vdd sg13_lv_pmos w=3.6525u l=3.38u ng=4 m=1
XM9 iout iout vdd vdd sg13_lv_pmos w=3.6525u l=3.38u ng=4 m=1
XC1 net3 vout cap_cmim w=9.98e-6 l=7.7e-6 m=4
XM6 vout net3 vss vss sg13_lv_nmos w=2.28u l=9.75u ng=1 m=1
**.ends
.end
