** sch_path: /home/pedersen/projects/IHP-AnalogAcademy/modules/module_1_bandgap_reference/part_3_layout/OTA_layout/full_OTA/schematic_mod/two_stage_OTA_layout.sch
.subckt two_stage_OTA_layout v- v+ vss vdd iout vout
*.PININFO v-:B v+:B vss:B vdd:B iout:B vout:B
M1 dn3 v- dn2 bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M2 dn4 v+ dn2 bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M8 dn4 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M10 dn3 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M15 dn2 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
M16 dn2 vdd vdd bulk sg13_lv_pmos l=3.7u w=3.64u ng=1 m=2
R1 vdd bulk ntap1 A = 0.1979378e-9 P = 0.243602e-3
M7 dn2 iout vdd bulk1 sg13_lv_pmos l=1.95u w=5.3u ng=1 m=1
R2 vss bulk2 ptap1 A = 15.54345e-12 P=53.44e-6
R3 vdd bulk1 ntap1 w=0.78e-6 l=0.78e-6
M3 dn3 dn3 vss bulk2 sg13_lv_nmos l=9.75u w=720n ng=1 m=1
M4 dn4 dn3 vss bulk2 sg13_lv_nmos l=9.75u w=720n ng=1 m=1
M5 vout iout vdd bulk4 sg13_lv_pmos l=2.08u w=75u ng=8 m=1
M6 vout dn4 vss bulk3 sg13_lv_nmos l=9.75u w=28.8u ng=4 m=1
M9 iout iout vdd bulk4 sg13_lv_pmos l=2.08u w=75u ng=8 m=1
C2 dn4 vout cap_cmim w=22.295e-6 l=22.295e-6 m=1
R4 vss bulk2 ptap1 A = 9.64655e-12, P = 0.18e-3
R5 vdd bulk3 ntap1 A = 27.435e-12, P = 0.177e-3
.ends
.end
