* Extracted by KLayout with SG13G2 LVS runset on : 27/03/2025 15:48

.SUBCKT input_common_centroid vdd dn3 v+ dn4 v\x2d
M$1 vdd vdd \$9 \$2 sg13_lv_pmos L=3.7u W=14.56u AS=4.9504p AD=4.9504p
+ PS=31.84u PD=31.84u
M$3 \$9 v+ dn4 \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p PS=15.92u
+ PD=15.92u
M$4 \$9 v\x2d dn3 \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p
+ PS=15.92u PD=15.92u
M$5 dn4 vdd vdd \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p PS=15.92u
+ PD=15.92u
M$6 dn3 vdd vdd \$2 sg13_lv_pmos L=3.7u W=7.28u AS=2.4752p AD=2.4752p PS=15.92u
+ PD=15.92u
R$13 \$2 vdd ntap1 A=28.7556p P=185.52u
.ENDS input_common_centroid
