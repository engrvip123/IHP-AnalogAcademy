* Extracted by KLayout with SG13G2 LVS runset on : 27/03/2025 16:03

.SUBCKT input_stage vss dn4 dn3 vdd dn2 iout
M$1 vss dn3 dn4 \$1 sg13_lv_nmos L=9.75u W=0.72u AS=0.2448p AD=0.2448p PS=2.12u
+ PD=2.12u
M$2 vss dn3 dn3 \$1 sg13_lv_nmos L=9.75u W=0.72u AS=0.2448p AD=0.2448p PS=2.12u
+ PD=2.12u
M$3 dn2 iout vdd \$8 sg13_lv_pmos L=1.95u W=5.3u AS=1.802p AD=1.802p PS=11.28u
+ PD=11.28u
R$4 \$8 vdd ntap1 A=7.5826p P=48.92u
R$5 \$1 vss ptap1 A=7.0975p P=56.78u
.ENDS input_stage
