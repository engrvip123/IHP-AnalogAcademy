** OTA_SIMPLE flat netlist
*.PININFO V-:B V+:B VSS:B VDD:B IOUT:B VOUT:B
M4 NET3 NET1 VSS VSS SG13_LV_NMOS L=9.75U W=720N NG=1 M=1
M3 NET1 NET1 VSS VSS SG13_LV_NMOS L=9.75U W=720N NG=1 M=1
M1 NET1 V- NET2 VDD SG13_LV_PMOS L=3.64U W=7.41U NG=1 M=1
M2 NET3 V+ NET2 VDD SG13_LV_PMOS L=3.64U W=7.41U NG=1 M=1
M5 NET2 IOUT VDD VDD SG13_LV_PMOS L=1.95U W=5.3U NG=1 M=1
M7 VOUT IOUT VDD VDD SG13_LV_PMOS L=2.08U W=75U NG=8 M=1
M6 VOUT NET3 VSS VSS SG13_LV_NMOS L=9.75U W=28.8U NG=4 M=1
M9 IOUT IOUT VDD VDD SG13_LV_PMOS L=2.08U W=75U NG=8 M=1
C2 NET3 VOUT CAP_CMIM W=22.295E-6 L=22.295E-6 M=1
.end
